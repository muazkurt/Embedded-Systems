library verilog;
use verilog.vl_types.all;
entity Status_Test is
end Status_Test;
